`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/03/12 14:53:28
// Design Name: 
// Module Name: MULT
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MULT(
    input clk,
    input reset,
    input [31:0] a,
    input [31:0] b,
    output [63:0] z
    );
    reg [31:0] ab00;
    reg [31:0] ab01;
    reg [31:0] ab02;
    reg [31:0] ab03;
    reg [31:0] ab04;
    reg [31:0] ab05;
    reg [31:0] ab06;
    reg [31:0] ab07;
    reg [31:0] ab08;
    reg [31:0] ab09;
    reg [31:0] ab10;
    reg [31:0] ab11;
    reg [31:0] ab12;
    reg [31:0] ab13;
    reg [31:0] ab14;
    reg [31:0] ab15;
    reg [31:0] ab16;
    reg [31:0] ab17;
    reg [31:0] ab18;
    reg [31:0] ab19;
    reg [31:0] ab20;
    reg [31:0] ab21;
    reg [31:0] ab22;
    reg [31:0] ab23;
    reg [31:0] ab24;
    reg [31:0] ab25;
    reg [31:0] ab26;
    reg [31:0] ab27;
    reg [31:0] ab28;
    reg [31:0] ab29;
    reg [31:0] ab30;
    reg [31:0] ab31;
    reg [63:0] temp;
    
    always @(posedge clk or negedge reset)
    begin
    if(reset)
    begin
        ab00<=0;
        ab01<=0;
        ab02<=0;
        ab03<=0;
        ab04<=0;
        ab05<=0;
        ab06<=0;
        ab07<=0;
        ab08<=0;
        ab09<=0;
        ab10<=0;
        ab11<=0;
        ab12<=0;
        ab13<=0;
        ab14<=0;
        ab15<=0;
        ab16<=0;
        ab17<=0;
        ab18<=0;
        ab19<=0;
        ab20<=0;
        ab21<=0;
        ab22<=0;
        ab23<=0;
        ab24<=0;
        ab25<=0;
        ab26<=0;
        ab27<=0;
        ab28<=0;
        ab29<=0;
        ab30<=0;
        ab31<=0;
        temp<=0;
    end
    else
    begin
        ab00<=b[0]?a:32'b0;
        ab01<=b[1]?a:32'b0;
        ab02<=b[2]?a:32'b0;
        ab03<=b[3]?a:32'b0;
        ab04<=b[4]?a:32'b0;
        ab05<=b[5]?a:32'b0;
        ab06<=b[6]?a:32'b0;
        ab07<=b[7]?a:32'b0;
        ab08<=b[8]?a:32'b0;
        ab09<=b[9]?a:32'b0;
        ab10<=b[10]?a:32'b0;
        ab11<=b[11]?a:32'b0;
        ab12<=b[12]?a:32'b0;
        ab13<=b[13]?a:32'b0;
        ab14<=b[14]?a:32'b0;
        ab15<=b[15]?a:32'b0;
        ab16<=b[16]?a:32'b0;
        ab17<=b[17]?a:32'b0;
        ab18<=b[18]?a:32'b0;
        ab19<=b[19]?a:32'b0;
        ab20<=b[20]?a:32'b0;
        ab21<=b[21]?a:32'b0;
        ab22<=b[22]?a:32'b0;
        ab23<=b[23]?a:32'b0;
        ab24<=b[24]?a:32'b0;
        ab25<=b[25]?a:32'b0;
        ab26<=b[26]?a:32'b0;
        ab27<=b[27]?a:32'b0;
        ab28<=b[28]?a:32'b0;
        ab29<=b[29]?a:32'b0;
        ab30<=b[30]?a:32'b0;
        ab31<=b[31]?a:32'b0;
    
       temp<=(({32'b1,~ab00[31],ab00[30:0]}        +
               {31'b0,~ab01[31],ab01[30:0], 1'b0}) +
              ({30'b0,~ab02[31],ab02[30:0], 2'b0}  +
               {29'b0,~ab03[31],ab03[30:0], 3'b0}))+
             (({28'b0,~ab04[31],ab04[30:0], 4'b0}  +
               {27'b0,~ab05[31],ab05[30:0], 5'b0}) +
              ({26'b0,~ab06[31],ab06[30:0], 6'b0}  +
               {25'b0,~ab07[31],ab07[30:0], 7'b0}))+
             (({24'b0,~ab08[31],ab08[30:0], 8'b0}  +
               {23'b0,~ab09[31],ab09[30:0], 9'b0}) +
              ({22'b0,~ab10[31],ab10[30:0],10'b0}  +
               {21'b0,~ab11[31],ab11[30:0],11'b0}))+
             (({20'b0,~ab12[31],ab12[30:0],12'b0}  +
               {19'b0,~ab13[31],ab13[30:0],13'b0}) +
              ({18'b0,~ab14[31],ab14[30:0],14'b0}  +
               {17'b0,~ab15[31],ab15[30:0],15'b0}))+
             (({16'b0,~ab16[31],ab16[30:0],16'b0}  +
               {15'b0,~ab17[31],ab17[30:0],17'b0}) +
              ({14'b0,~ab18[31],ab18[30:0],18'b0}  +
               {13'b0,~ab19[31],ab19[30:0],19'b0}))+
             (({12'b0,~ab20[31],ab20[30:0],20'b0}  +
               {11'b0,~ab21[31],ab21[30:0],21'b0}) +
              ({10'b0,~ab22[31],ab22[30:0],22'b0}  +
               { 9'b0,~ab23[31],ab23[30:0],23'b0}))+
             (({ 8'b0,~ab24[31],ab24[30:0],24'b0}  +
               { 7'b0,~ab25[31],ab25[30:0],25'b0}) +
              ({ 6'b0,~ab26[31],ab26[30:0],26'b0}  +
               { 5'b0,~ab27[31],ab27[30:0],27'b0}))+
             (({ 4'b0,~ab28[31],ab28[30:0],28'b0}  +
               { 3'b0,~ab29[31],ab29[30:0],29'b0}) +
              ({ 2'b0,~ab30[31],ab30[30:0],30'b0}  +
               { 1'b1,ab31[31],~ab31[30:0],31'b0}));
    end
    end
    assign z=temp;
endmodule
